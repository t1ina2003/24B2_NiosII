
module niosii (
	clk_clk,
	pio_led_export,
	pio_rst_export);	

	input		clk_clk;
	output	[7:0]	pio_led_export;
	input		pio_rst_export;
endmodule
